`timescale 1ns / 1ps 


module behavior_model_tb():
    reg[3:0] t_input; 
    wire t_F;
    integer i; 

